`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////

// fixed by using the correct syntax for assigning a value to a wire

//////////////////////////////////////////////////////////////////////////////////

module module3 (
    input  wire a,
    output wire b
);

  assign b = a;

endmodule
