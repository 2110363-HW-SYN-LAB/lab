`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////

// fixed by using the correct syntax for assigning a value to a reg

//////////////////////////////////////////////////////////////////////////////////

module module2 (
    input  wire a,
    output reg  b
);

  always @(*) begin
    b = a;
  end

endmodule
