`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////

// Fixed by correcting the syntax

//////////////////////////////////////////////////////////////////////////////////

module module1 (
    input  wire a,
    output wire b
);

assign b = a;

endmodule
