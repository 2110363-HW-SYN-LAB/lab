`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////

// This faulty module showcases an error message
// The error is cause by syntax error

//////////////////////////////////////////////////////////////////////////////////

module module1 (
    input  wire a,
    output wire b
);

assign 

endmodule
