`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////

// fixed by only driving the output wire with one input wire

//////////////////////////////////////////////////////////////////////////////////

module module4 (
    input  wire a,
    input  wire b,
    output wire c
);

  assign c = a & b;

endmodule
