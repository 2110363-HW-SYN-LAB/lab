`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////

// This faulty module showcases an error message
// The error is cause by using assign on reg

//////////////////////////////////////////////////////////////////////////////////

module module2 (
    input  wire a,
    output reg  b
);

  assign b = a;

endmodule
